�� sr Lesson_31.Student��-��˦  I ageL 	firstnamet Ljava/lang/String;L lastnameq ~ xp   t Mikhailt 	Belozerov